`ifndef MACROS_H_
`define MACROS_H_
typedef enum{transmit,recieve}  transaction;

`endif